`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:16:59 03/24/2021 
// Design Name: 
// Module Name:    Control_Unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Control_Unit(
    input[1:0] OpCode,
    output reg ALU_OP,
    output reg Reg_Write
    );
	
	always@(OpCode)
	 begin
		case(OpCode)
		2'b00: begin
						
						ALU_OP = 0; // Simple Addition
						Reg_Write = 1; // WriteBack is Needed
				 end
		2'b01: begin
						ALU_OP = 1; // Logical shift left
						Reg_Write = 1; // WriteBack is Needed
				 end
		default
				begin
						ALU_OP = 0; // Simple Addition
						Reg_Write = 0; // WriteBack is not Needed
				end
		endcase
	 end

endmodule
